module Notgate(
  input  wire in_,
  output wire out
);

  // Variables for output ports
  logic __out_bits;

  assign __out_bits = ~in_;

  assign out = __out_bits;
endmodule
